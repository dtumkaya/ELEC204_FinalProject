----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    14:45:44 06/07/2022 
-- Design Name: 
-- Module Name:    MinMaxMedianRange - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity MinMaxMedianRange is
    Port ( input1 : in  STD_LOGIC_VECTOR (3 downto 0);
           input2 : in  STD_LOGIC_VECTOR (3 downto 0);
           input3 : in  STD_LOGIC_VECTOR (3 downto 0);
           max : out  STD_LOGIC_VECTOR (3 downto 0);
           min : out  STD_LOGIC_VECTOR (3 downto 0);
           median : out  STD_LOGIC_VECTOR (3 downto 0);
           ranget : out  STD_LOGIC_VECTOR (3 downto 0));
end MinMaxMedianRange;

architecture Behavioral of MinMaxMedianRange is

begin


end Behavioral;

